VARNING!

'BF2MC Online' och 'BFMCSpy' definieras härmed som 'Tjänsterna' är fangjorda och drivna tjänster utformade för att återuppliva och bevara onlinefunktionerna i Battlefield 2: Modern Combat. Tjänsterna är inte på något sätt anslutna till eller drivs av EA, DICE, Gamespy eller närstående parter. All kontakt angående tjänsterna ska göras till vår Discord @ https://discord.gg/bf2mc.