   Välkommen till BF2:MC Online-tjänsten!

Genom att acceptera detta avtal samtycker du till följande spelserverregler och förstår att konsekvenserna av att bryta mot dessa regler kan resultera i att din åtkomst till servrarna återkallas eller att dina in-game-statistik justeras.

SPELSERVERREGLER:

Användning av alla tredjepartsverktyg för att få fördelar eller påverka spelupplevelsen är strängt förbjuden.

Användning av fusk för att få fördelar eller påverka spelupplevelsen är strängt förbjuden.

Alla former av glitchning för att få fördelar eller påverka spelupplevelsen är strängt förbjudna.

Misshandla eller trakassera inte andra spelare i spelet, såsom att medvetet teamdöda eller använda verbalt våld via din mikrofon.

Försök inte att utge dig för att vara andra medlemmar eller klaner inom gemenskapen eller tidigare spelare i spelet.

Missbruka inte funktionen för omröstningskick (votekick) i spelet.

Missbruka inte funktionen för in-game-meddelanden eller spelinbjudningar.

Missbruka inte spelets mekanik eller servrar för att manipulera de in-game-ledartavlorna (till exempel boosting eller padding).

Var inte inaktiv under långa perioder som skulle påverka spelupplevelsen.

Använd Mod Mail-boten på Discord för att rapportera regelbrytare.

Ha det så trevligt!

BFMCspy Team

discord.gg/bf2mc