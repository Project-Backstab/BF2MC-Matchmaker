Välkommen till BF2:MC Online Service!

Genom att acceptera detta avtal godkänner du följande spelserverregler och förstår att konsekvenserna av att bryta mot dessa regler kan resultera i att din åtkomst till servrarna återkallas.

SPELSERVER REGLER:

1. Användning av verktyg från tredje part för att få en fördel i spelet är strängt förbjudet.

2. All användning av fusk för att få en fördel i spelet är strängt förbjudet.

3. Alla former av glitching för att få en fördel är strängt förbjudna.

4. Missbruka eller trakassera inte andra spelare i spelet, såsom Målmedvetet Teamkilling och Verbal Abuse med din mikrofon.

5. Missbruka inte Votekick-funktionen i spelet.

6. Var en lagspelare och spela målet!

Använd [#report-a-player]-kanalen i discorden för att rapportera regelbrytare.


Var god njut!

Omega

discord.gg/bf2mc