   Välkommen till BFMCSpy!

När du skapar ett konto på vår tjänst, rekommenderas det starkt att du använder minnesvärda kontodetaljer. Det finns ingen "återställ lösenord" eller "återställ konto"-funktion tillgänglig för närvarande. Du kommer att kunna använda dessa uppgifter för att logga in på vår webbplats.

Genom att skapa och använda BFMCSpy-tjänsten godkänner du följande regler:

1. Utge dig inte som andra spelare
2. Inga kontonamn eller klannamn som innehåller förtal
3. Trakassera eller trakassera inte någon spelare när du skickar meddelanden
4. Håll Clan Motto's fria från förtal.

AVTAL:
DENNA PROGRAM TILLHANDAHÅLLS AV BIDRAGARE "I BEFINTLIGT SKICK" OCH NÅGON UTTRYCKLIG ELLER
UNDERFÖRSTÅDDA GARANTIER, INKLUSIVE, MEN INTE BEGRÄNSADE TILL, UNDERFÖRSTÅDDA GARANTIER OM SÄLJBARHET OCH LÄMPLIGHET FÖR ETT SÄRSKILT ÄNDAMÅL FRÅSES. UNDER INGA OMSTÄNDIGHETER SKA UPPHOVSRÄTTSINNEHAVAREN ELLER BIDRAGSGIVARNA VARA ANSVARIGA FÖR NÅGON DIREKTA, INDIREKTA, OAVSIKTLIGA, SPECIELLA, EXEMPELSKADOR ELLER FÖLJDSKADOR (INKLUSIVE, MEN INTE BEGRÄNSADE TILL, UPPHANDLING AV ERSÄTTNINGSSJÄNSTVAROR ELLER ERSÄTTNINGSSERVICE AV VAROR; .) OAVSETT ORSAKET OCH PÅ NÅGON TEORI OM ANSVAR, OAVSETT I KONTRAKT, STIKT ANSVAR ELLER SKADESTÅND (INKLUSIVE FÖRSIKTIGHET ELLER ANNAT SÄTT) SOM UPPSTÅR PÅ NÅGOT SÄTT UR ANVÄNDNING AV DENNA PROGRAM, ÄVEN OM DET HAR ORDET OM DET ÄR DET.